module mymultiplier(input [9:0] dataa, datab, output [19:0] w);
    assign w = dataa * datab;
endmodule